interface gen_cov_if();
  logic [7:0] A;
  logic [7:0] B;
  real curr_cov;
  
endinterface

