package my_pkg;
`include "Driver.sv"
`include "transaction.sv"
`include "generator.sv"
`include "Monitor.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "env.sv"
`include "Test.sv"
`include "functional_Coverage.sv"
`include "coverage_sub.sv"
//`include "rtl/alu.v"
endpackage
