package my_pkg;
`include "Driver.sv"
`include "Transaction.sv"
`include "generator.sv"
//`include "monitor.sv"
//`include "scoreboard.sv"
//`include "environment.SystemVerilog"
endpackage
