program automatic demo;
initial begin
$display("demo file");
end
endprogram
